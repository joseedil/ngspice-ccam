* CNTFET transfer curve
*
* To run, call ngspice with the -b option and use the spice_readfile.m
* Octave function.

*** Circuit description
* CNTFET
M1 vds vgs 0 0 mod1

* Voltage sources
V1 vgs 0 0.4
V2 vds 0 1

* CNTFET model
.MODEL mod1 nmos level=99
+idstn="0.25592" vthin="-0.17594" vth0in="35.662" athin="18.029"
+sthin="0.2" idstp="0" vthip="-0.032389" vth0ip="84.762" athip="9.0461"
+sthip="0.2" vdcr="1.5854" betdcr="1.0266" smss="10" facss="1"
+rscs="27.1845" rdcs="12.1844" ctn0="1.0274e-13" ctp0="1.0274e-13"
+vthqs="-0.1" vth0qs="0.66693" athqs="3" vthqd="-1.1" vth0qd="3.0386"
+athqd="2.6667" pqsd="0.16667" rmta="132236.5698" amto="117945.2195"
+cmt="1.8152e-17" pqmt="0.49425" rscm="47306.2244" rdcm="47306.2244"
+fanof="1" fanofmt="1" hoogef="0.002" beta_fn="1" rsf="0.001" rdf="0.001"
+rg="1" cgspar1="0" cgspar2="2.4844e-14" cgdpar1="2.7819e-15"
+cgdpar2="2.7819e-15" cdspar="2.4e-14" tnom="26.85" rths="0" rthm="0"
+zetrmta="0" zetamto="0" alvthin="0" alvth0in="0" alvthip="0" alvth0ip="0"
+alidst="0" alct0="0" alvthqs="0" alvth0qs="0" alvthqd="0" alvth0qd="0"
+alrscon="0" alrmcon="0" atrap="0" btrap="0" ctrap="0" w0trap="0" strap="0"


*** Analysis
* Just call ngspice -b cntfet.cir.
* It will simulate the circuit and output data on a file called rawspice.raw.

.control
dc V2 0 1 0.005 v1 0 1 0.1


* The following commands create a dump file with the data.
* To plot, call gnuplot and use the command
* gnuplot> plot "rawspice.raw" using 1:2

set wr_vecnames
set wr_singlescale
wrdata rawspice.raw -v2#branch vgs


* Alternative export command: more info exported.
*set filetype=ascii
*write rawspice.raw -v2#branch

.endc

.end
